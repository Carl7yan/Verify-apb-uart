interface clk_rst_interface (
    output logic reset_n,
    output logic clk
  );
  //import clk_rst_pkg::*;
endinterface
